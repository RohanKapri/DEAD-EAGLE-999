module main
fn period(planet string) f64 {
	return 31557600 * match planet {
		'Mercury' { 0.2408467 }
		'Venus' { 0.61519726 }
		'Earth' { 1.0 }
		'Mars' { 1.8808158 }
		'Jupiter' { 11.862615 }
		'Saturn' { 29.447498 }
		'Uranus' { 84.016846 }
		'Neptune' { 164.79132 }
		else { 0.0 }
	}
} 
fn age(seconds f64, planet string) !f64 {
	p := period(planet)
	if p == 0 {
		return error('${planet} is not a valid planet')
	}
	return seconds / p
}