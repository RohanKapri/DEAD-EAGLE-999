module main

fn truncate(phrase string) string {

  return phrase.limit(5)
}